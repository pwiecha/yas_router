// -------------------------------------------------------------
// Module: config_regs.v
// Author: PWI
// Release: 1.0, Jan 2019
// -------------------------------------------------------------

module config_regs (
  input [1:0] config_addr,
  input [1:0] config_data,
  input       config_en,
  output      ch0_addr,
  output      ch1_addr,
  output      ch2_addr,
  output      crc_en
);



endmodule
